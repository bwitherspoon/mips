`timescale 1ns / 1ps

module cpu_tb;

    localparam MEM_SIZE = 1024;
    localparam REG_SIZE = 32;
    localparam CLOCK_PERIOD = 10; // 100 MHz

    integer i;

    reg clk = 1;
    reg rst;

    cpu cpu (
        .clk(clk),
        .rst(rst)
    );

    always #(CLOCK_PERIOD/2) clk <= ~clk;

    initial begin
        $dumpfile("cpu.vcd");
        $dumpvars(1, cpu.clk, cpu.rst);
        $dumpvars(1, cpu.pc_if_id, cpu.ir_if_id);
        for (i = 0; i < MEM_SIZE; i = i + 1)
            $dumpvars(1, cpu.memory.mem_[i]);
        for (i = 0; i < REG_SIZE; i = i + 1)
            $dumpvars(1, cpu.regfile.regs_[i]);

        rst = 1;
        #(CLOCK_PERIOD+1) rst = 0;
        #(16*CLOCK_PERIOD);

        $display("All tests succeeded.");
        $finish;
    end

endmodule

